`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    03:42:08 03/06/2018 
// Design Name: 
// Module Name:    IM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module IM(PCout,Instruction_Out);
		input [63:0] PCout;
		output [31:0] Instruction_Out;
		reg [7:0] IM [0:255];
		
		initial 
		begin
		
		// LDUR X1, [X31, #8]
		// 11111000010_000001000_00_11111_00001
		IM[0] = 8'hF8;
		IM[1] = 8'h40;
		IM[2] = 8'h83;
		IM[3] = 8'hE1;
		
		//LDUR X2, [X31,#16]
		// 11111000010_000010000_00_11111_00010
		IM[4] = 8'hF8;
		IM[5] = 8'h41;
		IM[6] = 8'h03;
		IM[7] = 8'hE2;
		
		//LDUR X3, [X31,#24]
		// 11111000010_000011000_00_11111_00011
		IM[8] = 8'hF8;
		IM[9] = 8'h41;
		IM[10] = 8'h83;
		IM[11] = 8'hE3;
		
		//LDUR X4, [X31,#32]
		// 11111000010_000100000_00_11111_00100
		IM[12] = 8'hF8;
		IM[13] = 8'h42;
		IM[14] = 8'h03;
		IM[15] = 8'hE4;
		
		//LDUR X5, [X31,#40]
		// 11111000010_000101000_00_11111_00101
		IM[16] = 8'hF8;
		IM[17] = 8'h42;
		IM[18] = 8'h83;
		IM[19] = 8'hE5;
		
		//LDUR X6, [X31,#48]
		// 11111000010_000110000_00_11111_00110
		IM[20] = 8'hF8;
		IM[21] = 8'h43;
		IM[22] = 8'h03;
		IM[23] = 8'hE6;
		
		//LDUR X7, [X31,#56]
		// 11111000010_000111000_00_11111_00111
		IM[24] = 8'hF8;
		IM[25] = 8'h43;
		IM[26] = 8'h83;
		IM[27] = 8'hE7;
		
		
		//LDUR X8, [X31,#64]
		// 11111000010_001000000_00_11111_01000
		IM[28] = 8'hF8;
		IM[29] = 8'h44;
		IM[30] = 8'h03;
		IM[31] = 8'hE8;
		
		//LDUR X9, [X31,#72]
		// 11111000010_001001000_00_11111_01001
		IM[32] = 8'hF8;
		IM[33] = 8'h44;
		IM[34] = 8'h83;
		IM[35] = 8'hE9;
		
		
		//LDUR X10, [X31,#80]
		// 11111000010_001010000_00_11111_01010
		IM[36] = 8'hF8;
		IM[37] = 8'h45;
		IM[38] = 8'h03;
		IM[39] = 8'hEA;
		
		//LDUR X11, [X31,#88]
		// 11111000010_001011000_00_11111_01011
		IM[40] = 8'hF8;
		IM[41] = 8'h45;
		IM[42] = 8'h83;
		IM[43] = 8'hEB;
		
		//LDUR X12, [X31,#96]
		// 11111000010_001100000_00_11111_01100
		IM[44] = 8'hF8;
		IM[45] = 8'h46;
		IM[46] = 8'h03;
		IM[47] = 8'hEC;
		
		//ADD X2, X1, X3
		// 10001011000_00011_000000_00001_00010
		IM[48] = 8'h8B;
		IM[49] = 8'h03;
		IM[50] = 8'h00;
		IM[51] = 8'h22;
		
		
		//SUB X6, X5, X4
		// 11001011000_00100_000000_00101_00110
		IM[52] = 8'hCB;
		IM[53] = 8'h04;
		IM[54] = 8'h00;
		IM[55] = 8'hA6;
		
		//OR X9, X7, X8
		// 10101010000_01000_000000_00111_01001
		IM[56] = 8'hAA;
		IM[57] = 8'h08;
		IM[58] = 8'h00;
		IM[59] = 8'hE9; 
		
		
		//AND X12, X10, X11	
		// 10001010000_01011_000000_01010_01100
		IM[60] = 8'h8A;
		IM[61] = 8'h0B;
		IM[62] = 8'h01;
		IM[63] = 8'h4C; 
		
		
		end
		
		
		assign Instruction_Out = {IM[PCout+0],IM[PCout+1],IM[PCout+2],IM[PCout+3]};
		
		
endmodule
